`timescale 1ns/1ps
module led_sw(
    output led,
    input  sw
);

assign led = sw;

endmodule